// module moduleName #(
//     parameters
// ) (
//     ports
// );
    
// endmodule